module mips_cache_instr(
    input logic clk,
    input logic rst,
    
    input logic[31:0] addr,
    output logic[31:0] readdata,
    output logic stall
);



endmodule